library verilog;
use verilog.vl_types.all;
entity Adder4bit_tb is
end Adder4bit_tb;
